module test_DES3;
reg enc1_dec0;
reg [1:64] in, key;
wire [1:64] out;
			
	DES des (enc1_dec0, in, key, out);
	
	//Plain Text : 0000000000000001 -> 64'b1.
	//Key : 22234512987ABB23 -> 0010_0010_0010_0011_0100_0101_0001_0010_1001_1000_0111_1010_1011_1011_0010_0011.
	//Cypher Text : 0A4ED5C15A63FEA3 -> 0000_1010_0100_1110_1101_0101_1100_0001_0101_1010_0110_0011_1111_1110_1010_0011.

	initial begin 
		// Encrypting 
		enc1_dec0 = 1'b1;
		in = 64'b1;
		key = 64'b0010_0010_0010_0011_0100_0101_0001_0010_1001_1000_0111_1010_1011_1011_0010_0011;
		
		#100
		// Decrypting
		enc1_dec0 = 1'b0;
		in = out;
		key = 64'b0010_0010_0010_0011_0100_0101_0001_0010_1001_1000_0111_1010_1011_1011_0010_0011;
	end
		
endmodule
