module test_DES;
reg enc1_dec0;
reg [1:64] in, key;
wire [1:64] out;
			
	DES des (enc1_dec0, in, key, out);
	
	//Plain Text : 0123456789ABCDEF -> 0000_0001_0010_0011_0100_0101_0110_0111_1000_1001_1010_1011_1100_1101_1110_1111.
	//Key : 133457799BBCDFF1 -> 0001_0011_0011_0100_0101_0111_0111_1001_1001_1011_1011_1100_1101_1111_1111_0001.
	//Cypher Text : 85E813540F0AB405 -> 1000_0101_1110_1000_0001_0011_0101_0100_0000_1111_0000_1010_1011_0100_0000_0101.

	initial begin 
		// Encrypting 
		enc1_dec0 = 1'b1;
		in = 64'b0000_0001_0010_0011_0100_0101_0110_0111_1000_1001_1010_1011_1100_1101_1110_1111;
		key = 64'b0001_0011_0011_0100_0101_0111_0111_1001_1001_1011_1011_1100_1101_1111_1111_0001;
		
		#100
		// Decrypting
		enc1_dec0 = 1'b0;
		in = out;
		key = 64'b0001_0011_0011_0100_0101_0111_0111_1001_1001_1011_1011_1100_1101_1111_1111_0001;
	end
		
endmodule