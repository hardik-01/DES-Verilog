module test_DES2;
reg enc1_dec0;
reg [1:64] in, key;
wire [1:64] out;
			
	DES des (enc1_dec0, in, key, out);
	
	//Plain Text : 123456ABCD132536 -> 0001_0010_0011_0100_0101_0110_1010_1011_1100_1101_0001_0011_0010_0101_0011_0110.
	//Key : AABB09182736CCDD -> 1010_1010_1011_1011_0000_1001_0001_1000_0010_0111_0011_0110_1100_1100_1101_1101.
	//Cypher Text : C0B7A8D05F3A829C -> 1100_0000_1011_0111_1010_1000_1101_0000_0101_1111_0011_1010_1000_0010_1001_1100.

	initial begin 
		// Encrypting 
		enc1_dec0 = 1'b1;
		in = 64'b0001_0010_0011_0100_0101_0110_1010_1011_1100_1101_0001_0011_0010_0101_0011_0110;
		key = 64'b1010_1010_1011_1011_0000_1001_0001_1000_0010_0111_0011_0110_1100_1100_1101_1101;
		
		#100
		// Decrypting
		enc1_dec0 = 1'b0;
		in = out;
		key = 64'b1010_1010_1011_1011_0000_1001_0001_1000_0010_0111_0011_0110_1100_1100_1101_1101;
	end
		
endmodule
